module ROM0 (
    input logic [3:0] addRom,
    output logic [31:0] dataRom
);
    logic [31:0] rom [15:0];

    initial begin
        rom[0]  = 32'b00000000000000000000000000000000;
        rom[1]  = 32'b00000000000000000000000000000000;
        rom[2]  = 32'b00000000000000000000000000000000;
        rom[3]  = 32'b00000000000111111110000000000000;
        rom[4]  = 32'b00000000001111111111000000000000;
        rom[5]  = 32'b00000000000111111110000000000000;
        rom[6]  = 32'b00000000000000000000000000000000;
        rom[7]  = 32'b00000000000000000000000000000000;
        rom[8]  = 32'b00000000000000000000000000000000;
        rom[9]  = 32'b00000000000000000000000000000000;
        rom[10] = 32'b00000000000000000000000000000000;
        rom[11] = 32'b00000000000000000000000000000000;
        rom[12] = 32'b00000000000000000000000000000000;
        rom[13] = 32'b00000000000000000000000000000000;
        rom[14] = 32'b00000000000000000000000000000000;
        rom[15] = 32'b00000000000000000000000000000000;
    end

    assign dataRom = rom[addRom];
	 
endmodule
//.	

module ROM1 (
    input logic [3:0] addRom,
    output logic [31:0] dataRom
);
    logic [31:0] rom [15:0];

    initial begin
        rom[0]  = 32'b00000000000000000000000000000000;
        rom[1]  = 32'b00000000000000000000000000000000;
        rom[2]  = 32'b00000000000000000000000000000000;
        rom[3]  = 32'b00000000000111111110000000000000;
        rom[4]  = 32'b00000000001111111111000000000000;
        rom[5]  = 32'b00000000000111111110000000000000;
        rom[6]  = 32'b00000000000000000000000000000000;
        rom[7]  = 32'b00000000000000000000000000000000;
        rom[8]  = 32'b00000000000000000000000000000000;
        rom[9]  = 32'b00000000000000000000000000000000;
        rom[10] = 32'b00000000000000000000000000000000;
        rom[11] = 32'b00000000000000000000000000000000;
        rom[12] = 32'b00000000000000000000000000000000;
        rom[13] = 32'b00000000000000000000000000000000;
        rom[14] = 32'b00000000000000000000000000000000;
        rom[15] = 32'b00000000000000000000000000000000;
    end

    assign dataRom = rom[addRom];
endmodule


module ROM2 (
    input logic [3:0] addRom,
    output logic [31:0] dataRom
);
    logic [31:0] rom [15:0];

    initial begin
        rom[0]  = 32'b00000000000000000000000000000000;
        rom[1]  = 32'b00000000000000000000000000000000;
        rom[2]  = 32'b00000000000011111111000000000000;
        rom[3]  = 32'b00000000011111111111111000000000;
        rom[4]  = 32'b00000000111111111111111100000000;
        rom[5]  = 32'b00000000111111111111110000000000;
        rom[6]  = 32'b00000000001111111111000000000000;
        rom[7]  = 32'b01111111110011111111000000000000;
        rom[8]  = 32'b01111111111111111111000000000000;
        rom[9]  = 32'b00000111011111111110000000000000;
        rom[10] = 32'b00000000011110011110000000000000;
        rom[11] = 32'b00000000011110011110000000000000;
        rom[12] = 32'b00000000011110011110000000000000;
        rom[13] = 32'b00000000011110011110000000000000;
        rom[14] = 32'b00000011111100111111100000000000;
        rom[15] = 32'b00000000000000000000000000000000;
    end

    assign dataRom = rom[addRom];
endmodule


module ROM3 (
    input logic [3:0] addRom,
    output logic [31:0] dataRom
);
    logic [31:0] rom [15:0];

    initial begin
        rom[0]  = 32'b00000000000000000000000000000000;
        rom[1]  = 32'b00000000000000000000000000000000;
        rom[2]  = 32'b00000000000011111111000000000000;
        rom[3]  = 32'b00000000011111111111111000000000;
        rom[4]  = 32'b00000000111111111111111100000000;
        rom[5]  = 32'b00000000111111111111110000000000;
        rom[6]  = 32'b00000000001111111111000000000000;
        rom[7]  = 32'b00000000000011111111011111111100;
        rom[8]  = 32'b00000000011111111111111111111100;
        rom[9]  = 32'b00000000011111111110111100000000;
        rom[10] = 32'b00000000011110011110000000000000;
        rom[11] = 32'b00000000011110011110000000000000;
        rom[12] = 32'b00000000011110011110000000000000;
        rom[13] = 32'b00000000011110011110000000000000;
        rom[14] = 32'b00000011111100111111100000000000;
        rom[15] = 32'b00000000000000000000000000000000;
    end

    assign dataRom = rom[addRom];
endmodule
